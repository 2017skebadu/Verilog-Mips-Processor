// Module: instmem
// Description: instruction memory containing test program code.
// 
//

module instmem(
	input [31:0] pc,
	output [31:0] instOut
	);

reg [31:0] RAM [0:64] = {
	32'h20100001,
	32'h00102020,
	32'h0c00000a,
	32'h02108820,
	32'h00112020,
	32'h0c00000a,
	32'h02308020,
	32'h00102020,
	32'h0c00000a,
	32'h08000003,
	32'h30880001,
	32'h20020000,
	32'h15000001,
	32'h20020001,
	32'h03e00008,
	32'h0c000008,
	32'h21ce0001,
	32'had880000,
	32'h00000000,
	32'h00000000,
	32'h00000000,
	32'h00000000,
	32'h00000000,
	32'h00000000,
	32'h00000000,
	32'h00000000,
	32'h00000000,
	32'h00000000,
	32'h00000000,
	32'h00000000,
	32'h00000000,
	32'h00000000,
	32'h00000000,
	32'h00000000,
	32'h00000000,
	32'h00000000,
	32'h00000000,
	32'h00000000,
	32'h00000000,
	32'h00000000,
	32'h00000000,
	32'h00000000,
	32'h00000000,
	32'h00000000,
	32'h00000000,
	32'h00000000,
	32'h00000000,
	32'h00000000,
	32'h00000000,
	32'h00000000,
	32'h00000000,
	32'h00000000,
	32'h00000000,
	32'h00000000,
	32'h00000000,
	32'h00000000,
	32'h00000000,
	32'h00000000,
	32'h00000000,
	32'h00000000,
	32'h00000000,
	32'h00000000,
	32'h00000000,
	32'h00000000,
	32'h00000000
}; //must prefill memory with instruction code here when testing

assign instOut= RAM[int'(pc)];

endmodule
